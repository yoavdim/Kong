// HartsMatrixBitMap File
// A two level bitmap. dosplaying harts on the screen FWbruary  2021
// (c) Technion IIT, Department of Electrical Engineering 2021



module	winDraw	(
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position
					input logic	[10:0] offsetY,
					input logic activate,
					input logic on_enter,


					output	logic	drawingRequest, //output that the pixel should be dispalyed
					output	logic	[7:0] RGBout,  //rgb value from the bitmap
					output logic next_lvl
 ) ;


// Size represented as Number of X and Y bits
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 32*16 and use only the top left 20*15 pixels
// this is the bitmap  of the maze , if there is a one  the na whole 32*32 rectange will be drawn on the screen
// all numbers here are hard coded to simplify the  understanding


logic [0:14] [0:19]  MazeBiMapMask=
{
20'b	00000000000000000000, // win draw
20'b	10010010000000000000,
20'b	01010100000000000000,
20'b	00101000000000000000,
20'b	00000000000000000000,
20'b	00000000110000000000,
20'b	00000001001000000000,
20'b	00000001001000000000,
20'b	00000000110000000000,
20'b	00000000000000000000,
20'b	00000000000010010010,
20'b	00000000000001010100,
20'b	00000000000000101000,
20'b	00000000000000000000,
20'b	00000000000000000000
};


// pipeline (ff) to get the pixel color from the array
assign next_lvl = drawingRequest && on_enter;
//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		drawingRequest <= '0;
		//next_lvl <= '0;
	end
	else begin
		if (MazeBiMapMask[offsetY[9:5] ][offsetX[9:5]] == 1'b1 ) // take bits 5,6,7,8,9,10 from address to select  position in the maze
						RGBout <= 7'hd1 ;
		else
			RGBout <= 7'h3F;

		//next_lvl <= '0;
		if(activate )
			drawingRequest <= '1;
		if (on_enter) begin
			drawingRequest <= '0;
			//if(drawingRequest)
				//next_lvl <= '1;
		end


	end
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not
endmodule
